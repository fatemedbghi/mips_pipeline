module regFile(input clk, regWrite, input[4:0] readReg1,readReg2, writeReg, input[31:0] writeData, output reg[31:0] regData1,regData2,output equal);
  reg[0:31] regData[31:0];
  /*assign regData1 = (readReg1 == 5'b0)? 32'b0:regData[readReg1];*/
  always@(readReg1, regData[readReg1])begin
    if(readReg1 == 5'b0) regData1 <= 32'b0;
    else regData1 <= regData[readReg1];
  end
  /*assign regData2 = (readReg2 == 5'b0)? 32'b0:regData[readReg2];*/
  always@(readReg2, regData[readReg2])begin
    if(readReg2 == 5'b0) regData2 <= 32'b0;
    else regData2 <= regData[readReg2];
  end
  assign equal = (regData1 == regData2)?1'b1:1'b0;
  always@(negedge clk) begin
		if(regWrite) regData[writeReg] <= writeData;
	end
endmodule